module top_module (
    input  [31:0] in,
    output [31:0] out
);  //

  // assign out[31:24] = ...;

endmodule
